/*
    Module Name: stop_watch
    Description: Very simple stop watch
*/

module stop_watch (
    input logic clk, nRst_i,
    input logic button_i,
    output logic [2:0] mode_o,
    output logic [4:0] time_o
);
    // Write your code here!
endmodule